typedef uvm_sequencer#(sequence_item) ahb_seqr;