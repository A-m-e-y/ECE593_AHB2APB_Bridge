// This scoreboard validates the data flow between DUT and TB.
// Will be developed for MS5