// This scoreboard validates the data flow between DUT and TB.