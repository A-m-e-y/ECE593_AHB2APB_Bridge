// Coverage is now integrated into the scoreboard (scoreboard.sv)
// This file is kept for potential future standalone coverage extensions
