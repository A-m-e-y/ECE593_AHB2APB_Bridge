// Coverage is now integrated into the transaction class (txn.sv)
// This file is kept for potential future standalone coverage extensions
