// ============================================================================
// Comprehensive Coverage Module for AHB2APB Bridge
// ============================================================================
// This module provides extensive functional and code coverage including:
// - AHB Protocol Coverage
// - APB Protocol Coverage  
// - FSM State and Transition Coverage
// - Cross Coverage
// - CDC Coverage
// - Address Mapping Coverage
// ============================================================================

module coverage_collector(
    input wire Hclk,
    input wire Pclk,
    input wire Hresetn,
    
    // AHB Interface
    input wire [31:0] Haddr,
    input wire [31:0] Hwdata,
    input wire [31:0] Hrdata,
    input wire [1:0]  Htrans,
    input wire        Hwrite,
    input wire        Hreadyin,
    input wire        Hreadyout,
    input wire [1:0]  Hresp,
    input wire [2:0]  Hsize,
    input wire [2:0]  Hburst,
    
    // APB Interface
    input wire [31:0] Paddr,
    input wire [31:0] Pwdata,
    input wire [31:0] Prdata,
    input wire [2:0]  Pselx,
    input wire        Penable,
    input wire        Pwrite,
    
    // FSM State (from APB_FSM_Controller)
    input wire [2:0]  fsm_state,
    
    // Internal signals
    input wire        valid
);

// ============================================================================
// FSM State Definitions (match RTL)
// ============================================================================
typedef enum bit [2:0] {
    ST_IDLE     = 3'b000,
    ST_WWAIT    = 3'b001,
    ST_READ     = 3'b010,
    ST_WRITE    = 3'b011,
    ST_WRITEP   = 3'b100,
    ST_RENABLE  = 3'b101,
    ST_WENABLE  = 3'b110,
    ST_WENABLEP = 3'b111
} fsm_state_t;

// ============================================================================
// AHB Transaction Types
// ============================================================================
typedef enum bit [1:0] {
    IDLE   = 2'b00,
    BUSY   = 2'b01,
    NONSEQ = 2'b10,
    SEQ    = 2'b11
} htrans_type_t;

// ============================================================================
// 1. AHB PROTOCOL COVERAGE
// ============================================================================
covergroup cg_ahb_protocol @(posedge Hclk);
    option.per_instance = 1;
    option.name = "ahb_protocol_cov";
    
    // Basic AHB signals
    cp_hwrite: coverpoint Hwrite {
        bins read  = {0};
        bins write = {1};
    }
    
    cp_htrans: coverpoint Htrans {
        bins idle    = {IDLE};
        bins busy    = {BUSY};
        bins nonseq  = {NONSEQ};
        bins seq     = {SEQ};
    }
    
    cp_hsize: coverpoint Hsize {
        bins size_byte     = {3'b000};
        bins size_halfword = {3'b001};
        bins size_word     = {3'b010};
        bins size_dword    = {3'b011};
        bins size_line_4   = {3'b100};
        bins size_line_8   = {3'b101};
        bins others        = default;
    }
    
    cp_hburst: coverpoint Hburst {
        bins single = {3'b000};
        bins incr   = {3'b001};
        bins wrap4  = {3'b010};
        bins incr4  = {3'b011};
        bins wrap8  = {3'b100};
        bins incr8  = {3'b101};
        bins wrap16 = {3'b110};
        bins incr16 = {3'b111};
    }
    
    cp_hresp: coverpoint Hresp {
        bins okay  = {2'b00};
        bins error = {2'b01};
        bins retry = {2'b10};
        bins split = {2'b11};
    }
    
    // Cross coverage: Write/Read with different transfer types
    cx_write_trans: cross cp_hwrite, cp_htrans {
        ignore_bins idle_trans = binsof(cp_htrans) intersect {IDLE, BUSY};
    }
    
    // Cross coverage: Size with burst type
    cx_size_burst: cross cp_hsize, cp_hburst {
        ignore_bins invalid = binsof(cp_hsize) intersect {3'b100, 3'b101};
    }
    
    // Valid signal coverage
    cp_valid: coverpoint valid {
        bins asserted   = {1};
        bins deasserted = {0};
    }
    
    // Hreadyout coverage
    cp_hreadyout: coverpoint Hreadyout {
        bins ready    = {1};
        bins not_ready = {0};
    }
    
endgroup

// ============================================================================
// 2. APB PROTOCOL COVERAGE
// ============================================================================
covergroup cg_apb_protocol @(posedge Pclk);
    option.per_instance = 1;
    option.name = "apb_protocol_cov";
    
    // APB slave selection
    cp_pselx: coverpoint Pselx {
        bins slave0 = {3'b001};
        bins slave1 = {3'b010};
        bins slave2 = {3'b100};
        bins none   = {3'b000};
        bins invalid = default;
    }
    
    // APB enable
    cp_penable: coverpoint Penable {
        bins setup  = {0};
        bins access = {1};
    }
    
    // APB write/read
    cp_pwrite: coverpoint Pwrite {
        bins read  = {0};
        bins write = {1};
    }
    
    // APB Phase transitions (SETUP→ACCESS)
    cp_apb_phase: coverpoint {Pselx != 0, Penable} {
        bins setup_phase  = {2'b10};  // PSEL=1, PENABLE=0
        bins access_phase = {2'b11};  // PSEL=1, PENABLE=1
        bins idle_phase   = {2'b00};  // PSEL=0, PENABLE=0
    }
    
    // Cross: Slave selection with read/write
    cx_slave_rw: cross cp_pselx, cp_pwrite {
        ignore_bins no_slave = binsof(cp_pselx) intersect {3'b000};
    }
    
    // Cross: Slave selection with enable
    cx_slave_enable: cross cp_pselx, cp_penable {
        ignore_bins no_slave = binsof(cp_pselx) intersect {3'b000};
    }
    
endgroup

// ============================================================================
// 3. FSM STATE COVERAGE
// ============================================================================
covergroup cg_fsm_states @(posedge Hclk);
    option.per_instance = 1;
    option.name = "fsm_state_cov";
    
    // All FSM states
    cp_state: coverpoint fsm_state {
        bins idle     = {ST_IDLE};
        bins wwait    = {ST_WWAIT};
        bins read     = {ST_READ};
        bins write    = {ST_WRITE};
        bins writep   = {ST_WRITEP};
        bins renable  = {ST_RENABLE};
        bins wenable  = {ST_WENABLE};
        bins wenablep = {ST_WENABLEP};
    }
    
    // Cross: FSM state with valid signal
    cx_state_valid: cross cp_state, valid {
        bins idle_with_valid     = binsof(cp_state) intersect {ST_IDLE} && binsof(valid) intersect {1};
        bins idle_without_valid  = binsof(cp_state) intersect {ST_IDLE} && binsof(valid) intersect {0};
        bins wwait_with_valid    = binsof(cp_state) intersect {ST_WWAIT} && binsof(valid) intersect {1};
        bins wwait_without_valid = binsof(cp_state) intersect {ST_WWAIT} && binsof(valid) intersect {0};
    }
    
    // Cross: FSM state with Hreadyout
    cx_state_ready: cross cp_state, Hreadyout;
    
endgroup

// ============================================================================
// 4. FSM TRANSITION COVERAGE
// ============================================================================
covergroup cg_fsm_transitions @(posedge Hclk);
    option.per_instance = 1;
    option.name = "fsm_transition_cov";
    
    // State transitions
    cp_state_trans: coverpoint fsm_state {
        // All valid state transitions
        bins idle_to_wwait    = (ST_IDLE => ST_WWAIT);
        bins idle_to_read     = (ST_IDLE => ST_READ);
        bins idle_stay        = (ST_IDLE => ST_IDLE);
        
        bins wwait_to_write   = (ST_WWAIT => ST_WRITE);
        bins wwait_to_writep  = (ST_WWAIT => ST_WRITEP);
        
        bins read_to_renable  = (ST_READ => ST_RENABLE);
        
        bins write_to_wenable  = (ST_WRITE => ST_WENABLE);
        bins write_to_wenablep = (ST_WRITE => ST_WENABLEP);
        
        bins writep_to_wenablep = (ST_WRITEP => ST_WENABLEP);
        
        bins renable_to_idle  = (ST_RENABLE => ST_IDLE);
        bins renable_to_wwait = (ST_RENABLE => ST_WWAIT);
        bins renable_to_read  = (ST_RENABLE => ST_READ);
        
        bins wenable_to_idle  = (ST_WENABLE => ST_IDLE);
        bins wenable_to_wwait = (ST_WENABLE => ST_WWAIT);
        bins wenable_to_read  = (ST_WENABLE => ST_READ);
        
        bins wenablep_to_write  = (ST_WENABLEP => ST_WRITE);
        bins wenablep_to_writep = (ST_WENABLEP => ST_WRITEP);
        bins wenablep_to_read   = (ST_WENABLEP => ST_READ);
        
        // Sequences: Common transaction patterns
        bins write_sequence = (ST_IDLE => ST_WWAIT => ST_WRITE => ST_WENABLE => ST_IDLE);
        bins read_sequence  = (ST_IDLE => ST_READ => ST_RENABLE => ST_IDLE);
        bins pipelined_writes = (ST_IDLE => ST_WWAIT => ST_WRITEP => ST_WENABLEP => ST_WRITE => ST_WENABLE);
        bins write_then_read = (ST_WENABLE => ST_READ => ST_RENABLE => ST_IDLE);
        bins read_then_write = (ST_RENABLE => ST_WWAIT => ST_WRITE);
    }
    
endgroup

// ============================================================================
// 5. ADDRESS MAPPING COVERAGE
// ============================================================================
covergroup cg_address_mapping @(posedge Hclk iff (Htrans == NONSEQ || Htrans == SEQ));
    option.per_instance = 1;
    option.name = "address_mapping_cov";
    
    // AHB Address ranges for different APB slaves
    cp_haddr: coverpoint Haddr {
        bins slave0_range = {[32'h8000_0000 : 32'h83FF_FFFF]};  // Pselx[0]
        bins slave1_range = {[32'h8400_0000 : 32'h87FF_FFFF]};  // Pselx[1]
        bins slave2_range = {[32'h8800_0000 : 32'h8BFF_FFFF]};  // Pselx[2]
        bins other_range  = default;
    }
    
    // APB Address should match AHB address
    cp_paddr: coverpoint Paddr {
        bins slave0_range = {[32'h8000_0000 : 32'h83FF_FFFF]};
        bins slave1_range = {[32'h8400_0000 : 32'h87FF_FFFF]};
        bins slave2_range = {[32'h8800_0000 : 32'h8BFF_FFFF]};
        bins other_range  = default;
    }
    
    // Cross: Haddr with Pselx
    cx_addr_slave: cross cp_haddr, Pselx {
        bins slave0_addr = binsof(cp_haddr.slave0_range) && binsof(Pselx) intersect {3'b001};
        bins slave1_addr = binsof(cp_haddr.slave1_range) && binsof(Pselx) intersect {3'b010};
        bins slave2_addr = binsof(cp_haddr.slave2_range) && binsof(Pselx) intersect {3'b100};
    }
    
endgroup

// ============================================================================
// 6. CDC COVERAGE
// ============================================================================
covergroup cg_cdc @(posedge Pclk);
    option.per_instance = 1;
    option.name = "cdc_coverage";
    
    // Penable transitions in Pclk domain
    cp_penable_trans: coverpoint Penable {
        bins low_to_high = (0 => 1);
        bins high_to_low = (1 => 0);
        bins stay_high   = (1 => 1);
        bins stay_low    = (0 => 0);
    }
    
    // Pselx changes
    cp_pselx_change: coverpoint Pselx {
        bins none_to_slave0 = (3'b000 => 3'b001);
        bins none_to_slave1 = (3'b000 => 3'b010);
        bins none_to_slave2 = (3'b000 => 3'b100);
        bins slave_to_none  = ([3'b001:3'b100] => 3'b000);
        bins slave_change   = (3'b001 => 3'b010), (3'b010 => 3'b100), (3'b001 => 3'b100);
    }
    
    // Cross: Penable with Pwrite (detect READ/WRITE in APB domain)
    cx_penable_pwrite: cross cp_penable_trans, Pwrite;
    
endgroup

// ============================================================================
// 7. TRANSACTION SEQUENCE COVERAGE
// ============================================================================
covergroup cg_transaction_sequences @(posedge Hclk);
    option.per_instance = 1;
    option.name = "transaction_sequences_cov";
    
    // Back-to-back transactions
    cp_htrans_seq: coverpoint Htrans {
        bins nonseq_to_idle   = (NONSEQ => IDLE);
        bins nonseq_to_nonseq = (NONSEQ => NONSEQ);
        bins nonseq_to_seq    = (NONSEQ => SEQ);
        bins seq_to_seq       = (SEQ => SEQ);
        bins seq_to_idle      = (SEQ => IDLE);
        bins idle_to_nonseq   = (IDLE => NONSEQ);
    }
    
    // Write/Read sequences
    cp_rw_seq: coverpoint Hwrite {
        bins write_to_write = (1 => 1);
        bins write_to_read  = (1 => 0);
        bins read_to_write  = (0 => 1);
        bins read_to_read   = (0 => 0);
    }
    
    // Cross: Transaction type sequences with read/write
    cx_trans_rw_seq: cross cp_htrans_seq, cp_rw_seq;
    
endgroup

// ============================================================================
// 8. CORNER CASE COVERAGE
// ============================================================================
covergroup cg_corner_cases @(posedge Hclk);
    option.per_instance = 1;
    option.name = "corner_cases_cov";
    
    // Reset behavior
    cp_reset: coverpoint Hresetn {
        bins reset_active   = {0};
        bins reset_inactive = {1};
        bins reset_deassert = (0 => 1);
    }
    
    // Boundary addresses
    cp_addr_boundary: coverpoint Haddr {
        bins addr_min       = {32'h8000_0000};
        bins addr_max       = {32'h8BFF_FFFF};
        bins addr_slave0_max = {32'h83FF_FFFF};
        bins addr_slave1_min = {32'h8400_0000};
        bins addr_slave1_max = {32'h87FF_FFFF};
        bins addr_slave2_min = {32'h8800_0000};
        bins addr_mid        = {32'h8600_0000};
    }
    
    // Data patterns
    cp_wdata_pattern: coverpoint Hwdata {
        bins all_zeros  = {32'h0000_0000};
        bins all_ones   = {32'hFFFF_FFFF};
        bins alternating = {32'hAAAA_AAAA, 32'h5555_5555};
        bins walking_ones = {32'h0000_0001, 32'h0000_0002, 32'h0000_0004, 32'h0000_0008};
    }
    
endgroup

// ============================================================================
// COVERAGE INSTANTIATION
// ============================================================================
cg_ahb_protocol           ahb_cov;
cg_apb_protocol           apb_cov;
cg_fsm_states             fsm_state_cov;
cg_fsm_transitions        fsm_trans_cov;
cg_address_mapping        addr_map_cov;
cg_cdc                    cdc_cov;
cg_transaction_sequences  trans_seq_cov;
cg_corner_cases           corner_cov;

initial begin
    ahb_cov         = new();
    apb_cov         = new();
    fsm_state_cov   = new();
    fsm_trans_cov   = new();
    addr_map_cov    = new();
    cdc_cov         = new();
    trans_seq_cov   = new();
    corner_cov      = new();
end

// ============================================================================
// COVERAGE REPORTING
// ============================================================================
function void display_coverage();
    real ahb_coverage, apb_coverage, fsm_coverage, trans_coverage;
    real addr_coverage, cdc_coverage, seq_coverage, corner_coverage;
    real total_coverage;
    
    ahb_coverage    = ahb_cov.get_inst_coverage();
    apb_coverage    = apb_cov.get_inst_coverage();
    fsm_coverage    = fsm_state_cov.get_inst_coverage();
    trans_coverage  = fsm_trans_cov.get_inst_coverage();
    addr_coverage   = addr_map_cov.get_inst_coverage();
    cdc_coverage    = cdc_cov.get_inst_coverage();
    seq_coverage    = trans_seq_cov.get_inst_coverage();
    corner_coverage = corner_cov.get_inst_coverage();
    
    total_coverage = (ahb_coverage + apb_coverage + fsm_coverage + trans_coverage +
                      addr_coverage + cdc_coverage + seq_coverage + corner_coverage) / 8.0;
    
    $display("\n========== DETAILED COVERAGE REPORT ==========");
    $display("AHB Protocol Coverage:       %0.2f%%", ahb_coverage);
    $display("APB Protocol Coverage:       %0.2f%%", apb_coverage);
    $display("FSM State Coverage:          %0.2f%%", fsm_coverage);
    $display("FSM Transition Coverage:     %0.2f%%", trans_coverage);
    $display("Address Mapping Coverage:    %0.2f%%", addr_coverage);
    $display("CDC Coverage:                %0.2f%%", cdc_coverage);
    $display("Transaction Sequence Cov:    %0.2f%%", seq_coverage);
    $display("Corner Case Coverage:        %0.2f%%", corner_coverage);
    $display("----------------------------------------------");
    $display("TOTAL COVERAGE:              %0.2f%%", total_coverage);
    $display("==============================================\n");
endfunction

endmodule

